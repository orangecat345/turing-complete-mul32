module mul8_yjy (clk, rst, wi_a_8bit, wi_b_8bit, wo_compr1_16bit, wo_compr0_16bit);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [7:0] wi_a_8bit;
  input  wire [7:0] wi_b_8bit;
  output  wire [15:0] wo_compr1_16bit;
  output  wire [15:0] wo_compr0_16bit;

  TC_Splitter8 # (.UUID(64'd871884273925886032 ^ UUID)) Splitter8_0 (.in(wire_12), .out0(wire_55), .out1(wire_11), .out2(wire_108), .out3(wire_7), .out4(wire_71), .out5(wire_89), .out6(wire_62), .out7(wire_24));
  TC_Maker16 # (.UUID(64'd1141963268693816925 ^ UUID)) Maker16_1 (.in0(wire_21), .in1(8'd0), .out(wire_23));
  TC_Splitter16 # (.UUID(64'd1061786111241966781 ^ UUID)) Splitter16_2 (.in(wire_61), .out0(wire_21), .out1(wire_78));
  TC_Splitter16 # (.UUID(64'd4288354615799651112 ^ UUID)) Splitter16_3 (.in(wire_99), .out0(wire_13), .out1(wire_20));
  TC_Splitter8 # (.UUID(64'd3235360505789212136 ^ UUID)) Splitter8_4 (.in(wire_13), .out0(wire_57), .out1(wire_31), .out2(wire_80), .out3(wire_3), .out4(wire_28), .out5(wire_46), .out6(wire_9), .out7(wire_91));
  TC_Maker8 # (.UUID(64'd3412598782661834206 ^ UUID)) Maker8_5 (.in0(1'd0), .in1(1'd0), .in2(wire_57), .in3(wire_31), .in4(wire_80), .in5(wire_3), .in6(wire_28), .in7(wire_46), .out(wire_51));
  TC_Maker8 # (.UUID(64'd261245533796592106 ^ UUID)) Maker8_6 (.in0(wire_9), .in1(wire_91), .in2(1'd0), .in3(1'd0), .in4(1'd0), .in5(1'd0), .in6(1'd0), .in7(1'd0), .out(wire_84));
  TC_Maker16 # (.UUID(64'd1348990164601925966 ^ UUID)) Maker16_7 (.in0(wire_51), .in1(wire_84), .out(wire_26));
  TC_Splitter16 # (.UUID(64'd1739465113782735944 ^ UUID)) Splitter16_8 (.in(wire_22), .out0(wire_105), .out1(wire_16));
  TC_Splitter8 # (.UUID(64'd4192656587422330661 ^ UUID)) Splitter8_9 (.in(wire_105), .out0(wire_42), .out1(wire_39), .out2(wire_48), .out3(wire_59), .out4(wire_65), .out5(wire_5), .out6(wire_10), .out7(wire_107));
  TC_Maker8 # (.UUID(64'd3516508877784600463 ^ UUID)) Maker8_10 (.in0(1'd0), .in1(1'd0), .in2(1'd0), .in3(1'd0), .in4(wire_42), .in5(wire_39), .in6(wire_48), .in7(wire_59), .out(wire_34));
  TC_Maker16 # (.UUID(64'd3969345435572237875 ^ UUID)) Maker16_11 (.in0(wire_34), .in1(wire_85), .out(wire_53));
  TC_Maker8 # (.UUID(64'd3679138009761726937 ^ UUID)) Maker8_12 (.in0(wire_65), .in1(wire_5), .in2(wire_10), .in3(wire_107), .in4(1'd0), .in5(1'd0), .in6(1'd0), .in7(1'd0), .out(wire_85));
  TC_Splitter16 # (.UUID(64'd1657932571700045497 ^ UUID)) Splitter16_13 (.in(wire_18), .out0(wire_30), .out1(wire_66));
  TC_Maker8 # (.UUID(64'd842108616878208921 ^ UUID)) Maker8_14 (.in0(1'd0), .in1(1'd0), .in2(1'd0), .in3(1'd0), .in4(1'd0), .in5(1'd0), .in6(wire_104), .in7(wire_93), .out(wire_97));
  TC_Maker8 # (.UUID(64'd3628476313312055207 ^ UUID)) Maker8_15 (.in0(wire_19), .in1(wire_86), .in2(wire_88), .in3(wire_4), .in4(wire_64), .in5(wire_101), .in6(1'd0), .in7(1'd0), .out(wire_56));
  TC_Maker16 # (.UUID(64'd3537796938386562727 ^ UUID)) Maker16_16 (.in0(wire_97), .in1(wire_56), .out(wire_17));
  TC_Splitter8 # (.UUID(64'd3998799440510990507 ^ UUID)) Splitter8_17 (.in(wire_30), .out0(wire_104), .out1(wire_93), .out2(wire_19), .out3(wire_86), .out4(wire_88), .out5(wire_4), .out6(wire_64), .out7(wire_101));
  TC_Splitter16 # (.UUID(64'd2527945987833496148 ^ UUID)) Splitter16_18 (.in(wire_49), .out0(wire_43), .out1(wire_63));
  TC_Splitter8 # (.UUID(64'd1103205388868845716 ^ UUID)) Splitter8_19 (.in(wire_43), .out0(wire_67), .out1(wire_14), .out2(wire_27), .out3(wire_103), .out4(wire_41), .out5(wire_32), .out6(wire_50), .out7(wire_1));
  TC_Splitter8 # (.UUID(64'd1868573819058257977 ^ UUID)) Splitter8_20 (.in(wire_63), .out0(wire_102), .out1(wire_40), .out2(wire_25), .out3(wire_82), .out4(wire_70), .out5(wire_95), .out6(wire_72), .out7());
  TC_Maker8 # (.UUID(64'd3551920810937562814 ^ UUID)) Maker8_21 (.in0(1'd0), .in1(wire_67), .in2(wire_14), .in3(wire_27), .in4(wire_103), .in5(wire_41), .in6(wire_32), .in7(wire_50), .out(wire_100));
  TC_Maker8 # (.UUID(64'd2444816234400511777 ^ UUID)) Maker8_22 (.in0(wire_1), .in1(wire_102), .in2(wire_40), .in3(wire_25), .in4(wire_82), .in5(wire_70), .in6(wire_95), .in7(wire_72), .out(wire_58));
  TC_Maker16 # (.UUID(64'd1414549126463634680 ^ UUID)) Maker16_23 (.in0(wire_100), .in1(wire_58), .out(wire_36));
  TC_Splitter8 # (.UUID(64'd704655723420817405 ^ UUID)) Splitter8_24 (.in(wire_78), .out0(wire_44), .out1(wire_33), .out2(), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd1686439310734374058 ^ UUID)) Splitter8_25 (.in(wire_20), .out0(wire_98), .out1(wire_0), .out2(), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd3803561959248594564 ^ UUID)) Splitter8_26 (.in(wire_16), .out0(wire_37), .out1(wire_2), .out2(), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd3193712430592095588 ^ UUID)) Splitter8_27 (.in(wire_66), .out0(wire_75), .out1(wire_68), .out2(), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Maker8 # (.UUID(64'd4272259269328703660 ^ UUID)) Maker8_28 (.in0(wire_44), .in1(wire_33), .in2(wire_98), .in3(wire_0), .in4(wire_37), .in5(wire_2), .in6(wire_75), .in7(wire_68), .out(wire_79));
  TC_Maker16 # (.UUID(64'd15451527055606716 ^ UUID)) Maker16_29 (.in0(8'd0), .in1(wire_79), .out(wire_52));
  booth_10bit_yjy # (.UUID(64'd1813826030400042322 ^ UUID)) booth_10bit_yjy_30 (.clk(clk), .rst(rst), .wi_8_bit(wire_38), .wi_a_0(wire_55), .wi_a_1(wire_11), .wo_pp_10bit(wire_61));
  booth_10bit_yjy # (.UUID(64'd4016882924763955475 ^ UUID)) booth_10bit_yjy_31 (.clk(clk), .rst(rst), .wi_8_bit(wire_38), .wi_a_0(wire_108), .wi_a_1(wire_7), .wo_pp_10bit(wire_99));
  booth_10bit_yjy # (.UUID(64'd2315150674972468301 ^ UUID)) booth_10bit_yjy_32 (.clk(clk), .rst(rst), .wi_8_bit(wire_38), .wi_a_0(wire_71), .wi_a_1(wire_89), .wo_pp_10bit(wire_22));
  booth_10bit_yjy # (.UUID(64'd3870356565631179713 ^ UUID)) booth_10bit_yjy_33 (.clk(clk), .rst(rst), .wi_8_bit(wire_38), .wi_a_0(wire_62), .wi_a_1(wire_24), .wo_pp_10bit(wire_18));
  Compr42with16Bit_yjy # (.UUID(64'd2230197389688683817 ^ UUID)) Compr42with16Bit_yjy_34 (.clk(clk), .rst(rst), .Input_1(wire_23), .Input_2(wire_26), .Input_3(wire_53), .Input_4(wire_17), .Output_1(wire_49), .Output_2(wire_6));
  Compr42with16Bit_yjy # (.UUID(64'd3542027003057700292 ^ UUID)) Compr42with16Bit_yjy_35 (.clk(clk), .rst(rst), .Input_1(16'd0), .Input_2(wire_36), .Input_3(wire_6), .Input_4(wire_52), .Output_1(wire_47), .Output_2(wire_96));
  TC_Splitter8 # (.UUID(64'd2540382302098490914 ^ UUID)) Splitter8_36 (.in(wire_29), .out0(wire_87), .out1(wire_81), .out2(wire_8), .out3(wire_77), .out4(wire_54), .out5(wire_109), .out6(wire_15), .out7(wire_76));
  TC_Splitter8 # (.UUID(64'd1746776852373521768 ^ UUID)) Splitter8_37 (.in(wire_60), .out0(wire_45), .out1(wire_92), .out2(wire_73), .out3(wire_69), .out4(wire_94), .out5(wire_83), .out6(wire_35), .out7());
  TC_Splitter16 # (.UUID(64'd1318736299301609568 ^ UUID)) Splitter16_38 (.in(wire_47), .out0(wire_29), .out1(wire_60));
  TC_Maker8 # (.UUID(64'd4114772111335134137 ^ UUID)) Maker8_39 (.in0(1'd0), .in1(wire_87), .in2(wire_81), .in3(wire_8), .in4(wire_77), .in5(wire_54), .in6(wire_109), .in7(wire_15), .out(wire_106));
  TC_Maker8 # (.UUID(64'd327153469904015032 ^ UUID)) Maker8_40 (.in0(wire_76), .in1(wire_45), .in2(wire_92), .in3(wire_73), .in4(wire_69), .in5(wire_94), .in6(wire_83), .in7(wire_35), .out(wire_74));
  TC_Maker16 # (.UUID(64'd4515871205160287203 ^ UUID)) Maker16_41 (.in0(wire_106), .in1(wire_74), .out(wire_90));

  wire [0:0] wire_0;
  wire [0:0] wire_1;
  wire [0:0] wire_2;
  wire [0:0] wire_3;
  wire [0:0] wire_4;
  wire [0:0] wire_5;
  wire [15:0] wire_6;
  wire [0:0] wire_7;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  wire [0:0] wire_10;
  wire [0:0] wire_11;
  wire [7:0] wire_12;
  assign wire_12 = wi_b_8bit;
  wire [7:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  wire [7:0] wire_16;
  wire [15:0] wire_17;
  wire [15:0] wire_18;
  wire [0:0] wire_19;
  wire [7:0] wire_20;
  wire [7:0] wire_21;
  wire [15:0] wire_22;
  wire [15:0] wire_23;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  wire [15:0] wire_26;
  wire [0:0] wire_27;
  wire [0:0] wire_28;
  wire [7:0] wire_29;
  wire [7:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [7:0] wire_34;
  wire [0:0] wire_35;
  wire [15:0] wire_36;
  wire [0:0] wire_37;
  wire [7:0] wire_38;
  assign wire_38 = wi_a_8bit;
  wire [0:0] wire_39;
  wire [0:0] wire_40;
  wire [0:0] wire_41;
  wire [0:0] wire_42;
  wire [7:0] wire_43;
  wire [0:0] wire_44;
  wire [0:0] wire_45;
  wire [0:0] wire_46;
  wire [15:0] wire_47;
  wire [0:0] wire_48;
  wire [15:0] wire_49;
  wire [0:0] wire_50;
  wire [7:0] wire_51;
  wire [15:0] wire_52;
  wire [15:0] wire_53;
  wire [0:0] wire_54;
  wire [0:0] wire_55;
  wire [7:0] wire_56;
  wire [0:0] wire_57;
  wire [7:0] wire_58;
  wire [0:0] wire_59;
  wire [7:0] wire_60;
  wire [15:0] wire_61;
  wire [0:0] wire_62;
  wire [7:0] wire_63;
  wire [0:0] wire_64;
  wire [0:0] wire_65;
  wire [7:0] wire_66;
  wire [0:0] wire_67;
  wire [0:0] wire_68;
  wire [0:0] wire_69;
  wire [0:0] wire_70;
  wire [0:0] wire_71;
  wire [0:0] wire_72;
  wire [0:0] wire_73;
  wire [7:0] wire_74;
  wire [0:0] wire_75;
  wire [0:0] wire_76;
  wire [0:0] wire_77;
  wire [7:0] wire_78;
  wire [7:0] wire_79;
  wire [0:0] wire_80;
  wire [0:0] wire_81;
  wire [0:0] wire_82;
  wire [0:0] wire_83;
  wire [7:0] wire_84;
  wire [7:0] wire_85;
  wire [0:0] wire_86;
  wire [0:0] wire_87;
  wire [0:0] wire_88;
  wire [0:0] wire_89;
  wire [15:0] wire_90;
  assign wo_compr0_16bit = wire_90;
  wire [0:0] wire_91;
  wire [0:0] wire_92;
  wire [0:0] wire_93;
  wire [0:0] wire_94;
  wire [0:0] wire_95;
  wire [15:0] wire_96;
  assign wo_compr1_16bit = wire_96;
  wire [7:0] wire_97;
  wire [0:0] wire_98;
  wire [15:0] wire_99;
  wire [7:0] wire_100;
  wire [0:0] wire_101;
  wire [0:0] wire_102;
  wire [0:0] wire_103;
  wire [0:0] wire_104;
  wire [7:0] wire_105;
  wire [7:0] wire_106;
  wire [0:0] wire_107;
  wire [0:0] wire_108;
  wire [0:0] wire_109;

endmodule
