module mulMiddle_2_1_yjy (clk, rst, clk, rstn, Input, Output_1, Output_2);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [0:0] clk;
  input  wire [0:0] rstn;
  input  wire [63:0] Input;
  output  wire [7:0] Output_1;
  output  wire [15:0] Output_2;

  TC_Register # (.UUID(64'd2751721783843254026 ^ UUID), .BIT_WIDTH(64'd64)) Register64_0 (.clk(clk), .rst(rst), .load(wire_3), .save(wire_8), .in(wire_14), .out(wire_4));
  TC_Not # (.UUID(64'd579745791837774298 ^ UUID), .BIT_WIDTH(64'd1)) Not_1 (.in(wire_32), .out(wire_6));
  TC_Or # (.UUID(64'd416440449238657224 ^ UUID), .BIT_WIDTH(64'd1)) Or_2 (.in0(wire_23), .in1(wire_6), .out(wire_8));
  TC_Not # (.UUID(64'd1355564700480115559 ^ UUID), .BIT_WIDTH(64'd1)) Not_3 (.in(wire_8), .out(wire_3));
  TC_Mux # (.UUID(64'd3750024940026240015 ^ UUID), .BIT_WIDTH(64'd64)) Mux64_4 (.sel(wire_8), .in0(wire_4), .in1(wire_14), .out(wire_26));
  TC_Mux # (.UUID(64'd1729767011881167311 ^ UUID), .BIT_WIDTH(64'd64)) Mux64_5 (.sel(wire_6), .in0(wire_5), .in1(64'd0), .out(wire_14));
  TC_Splitter64 # (.UUID(64'd4323783475943063022 ^ UUID)) Splitter64_6 (.in(wire_26), .out0(wire_25), .out1(wire_31), .out2(wire_17), .out3(wire_16), .out4(wire_12), .out5(wire_24), .out6(wire_20), .out7(wire_27));
  TC_Maker32 # (.UUID(64'd1955231400302693653 ^ UUID)) Maker32_7 (.in0(wire_25), .in1(wire_31), .in2(wire_17), .in3(wire_16), .out(wire_2));
  TC_Maker32 # (.UUID(64'd2072935069226845658 ^ UUID)) Maker32_8 (.in0(wire_12), .in1(wire_24), .in2(wire_20), .in3(wire_27), .out(wire_19));
  TC_Splitter32 # (.UUID(64'd732592950980183219 ^ UUID)) Splitter32_9 (.in(wire_2), .out0(wire_22), .out1(wire_9), .out2(), .out3());
  TC_Splitter32 # (.UUID(64'd4244625817818765988 ^ UUID)) Splitter32_10 (.in(wire_19), .out0(wire_28), .out1(wire_13), .out2(), .out3());
  TC_Register # (.UUID(64'd849181173002087696 ^ UUID), .BIT_WIDTH(64'd16)) Register16_11 (.clk(clk), .rst(rst), .load(wire_3), .save(wire_8), .in(wire_21), .out(wire_18));
  TC_Mux # (.UUID(64'd1483690337929278922 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_12 (.sel(wire_6), .in0(wire_1), .in1(16'd0), .out(wire_21));
  TC_Register # (.UUID(64'd225614132390476503 ^ UUID), .BIT_WIDTH(64'd8)) Register8_13 (.clk(clk), .rst(rst), .load(wire_3), .save(wire_8), .in(wire_10), .out(wire_7));
  TC_Mux # (.UUID(64'd874535666843899459 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_14 (.sel(wire_6), .in0(wire_15), .in1(8'd0), .out(wire_10));
  TC_Mux # (.UUID(64'd3068677969550485877 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_15 (.sel(wire_8), .in0(wire_18), .in1(wire_21), .out(wire_11));
  TC_Mux # (.UUID(64'd1772225095273392886 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_16 (.sel(wire_8), .in0(wire_7), .in1(wire_10), .out(wire_29));
  mul8_top_yjy # (.UUID(64'd2797592024929963849 ^ UUID)) mul8_top_yjy_17 (.clk(clk), .rst(rst), .wi_a_8bit(wire_22), .wi_b_8bit(wire_13), .Output(wire_0));
  mul8_top_yjy # (.UUID(64'd2106126521548271831 ^ UUID)) mul8_top_yjy_18 (.clk(clk), .rst(rst), .wi_a_8bit(wire_9), .wi_b_8bit(wire_28), .Output(wire_30));
  adder_16bit_lgy # (.UUID(64'd2682928204690924665 ^ UUID)) adder_16bit_lgy_19 (.clk(clk), .rst(rst), .i_a_16(wire_0), .i_b_16(wire_30), .Cin(1'd0), .Output_1(wire_1), .Output_2(wire_15));

  wire [15:0] wire_0;
  wire [15:0] wire_1;
  wire [31:0] wire_2;
  wire [0:0] wire_3;
  wire [63:0] wire_4;
  wire [63:0] wire_5;
  assign wire_5 = Input;
  wire [0:0] wire_6;
  wire [7:0] wire_7;
  wire [0:0] wire_8;
  wire [7:0] wire_9;
  wire [7:0] wire_10;
  wire [15:0] wire_11;
  assign Output_2 = wire_11;
  wire [7:0] wire_12;
  wire [7:0] wire_13;
  wire [63:0] wire_14;
  wire [7:0] wire_15;
  wire [7:0] wire_16;
  wire [7:0] wire_17;
  wire [15:0] wire_18;
  wire [31:0] wire_19;
  wire [7:0] wire_20;
  wire [15:0] wire_21;
  wire [7:0] wire_22;
  wire [0:0] wire_23;
  assign wire_23 = clk;
  wire [7:0] wire_24;
  wire [7:0] wire_25;
  wire [63:0] wire_26;
  wire [7:0] wire_27;
  wire [7:0] wire_28;
  wire [7:0] wire_29;
  assign Output_1 = wire_29;
  wire [15:0] wire_30;
  wire [7:0] wire_31;
  wire [0:0] wire_32;
  assign wire_32 = rstn;

endmodule
