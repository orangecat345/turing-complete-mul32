module mulMiddle_4_1_yjy (clk, rst, clk, rstn, i_msg_64, Output_1, Output_2, Output_3);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [0:0] clk;
  input  wire [0:0] rstn;
  input  wire [63:0] i_msg_64;
  output  wire [7:0] Output_1;
  output  wire [7:0] Output_2;
  output  wire [7:0] Output_3;

  TC_Register # (.UUID(64'd1962039682932341795 ^ UUID), .BIT_WIDTH(64'd64)) Register64_0 (.clk(clk), .rst(rst), .load(wire_3), .save(wire_13), .in(wire_28), .out(wire_19));
  TC_Not # (.UUID(64'd1933006174712696322 ^ UUID), .BIT_WIDTH(64'd1)) Not_1 (.in(wire_63), .out(wire_2));
  TC_Or # (.UUID(64'd466796145083473585 ^ UUID), .BIT_WIDTH(64'd1)) Or_2 (.in0(wire_14), .in1(wire_2), .out(wire_13));
  TC_Not # (.UUID(64'd3042922256194320506 ^ UUID), .BIT_WIDTH(64'd1)) Not_3 (.in(wire_13), .out(wire_3));
  TC_Mux # (.UUID(64'd4575681795967979293 ^ UUID), .BIT_WIDTH(64'd64)) Mux64_4 (.sel(wire_2), .in0(wire_12), .in1(64'd0), .out(wire_28));
  TC_Mux # (.UUID(64'd3405608948629277411 ^ UUID), .BIT_WIDTH(64'd64)) Mux64_5 (.sel(wire_13), .in0(wire_19), .in1(wire_28), .out(wire_21));
  TC_Splitter64 # (.UUID(64'd2298753791118958783 ^ UUID)) Splitter64_6 (.in(wire_21), .out0(wire_61), .out1(wire_40), .out2(wire_9), .out3(wire_52), .out4(wire_57), .out5(wire_29), .out6(wire_33), .out7(wire_34));
  TC_Maker32 # (.UUID(64'd3976455095654061933 ^ UUID)) Maker32_7 (.in0(wire_61), .in1(wire_40), .in2(wire_9), .in3(wire_52), .out(wire_42));
  TC_Maker32 # (.UUID(64'd4001311498107799180 ^ UUID)) Maker32_8 (.in0(wire_57), .in1(wire_29), .in2(wire_33), .in3(wire_34), .out(wire_18));
  TC_Splitter32 # (.UUID(64'd1603467459090654200 ^ UUID)) Splitter32_9 (.in(wire_42), .out0(wire_50), .out1(wire_46), .out2(wire_60), .out3(wire_54));
  TC_Splitter32 # (.UUID(64'd4609873788031112092 ^ UUID)) Splitter32_10 (.in(wire_18), .out0(wire_64), .out1(wire_8), .out2(wire_59), .out3(wire_38));
  mul8_top_yjy # (.UUID(64'd1237322937714988485 ^ UUID)) mul8_top_yjy_11 (.clk(clk), .rst(rst), .wi_a_8bit(wire_50), .wi_b_8bit(wire_38), .Output(wire_53));
  mul8_top_yjy # (.UUID(64'd802669220327225322 ^ UUID)) mul8_top_yjy_12 (.clk(clk), .rst(rst), .wi_a_8bit(wire_46), .wi_b_8bit(wire_59), .Output(wire_44));
  mul8_top_yjy # (.UUID(64'd2960529241396483624 ^ UUID)) mul8_top_yjy_13 (.clk(clk), .rst(rst), .wi_a_8bit(wire_60), .wi_b_8bit(wire_8), .Output(wire_20));
  mul8_top_yjy # (.UUID(64'd3151330249751273606 ^ UUID)) mul8_top_yjy_14 (.clk(clk), .rst(rst), .wi_a_8bit(wire_54), .wi_b_8bit(wire_64), .Output(wire_0));
  Compr42with16Bits_yjy # (.UUID(64'd1284012806296956213 ^ UUID)) Compr42with16Bits_yjy_15 (.clk(clk), .rst(rst), .Input_1(wire_53), .Input_2(wire_44), .Input_3(wire_20), .Input_4(wire_0), .\1_out (wire_11), .sum(wire_17), .carr(wire_4));
  adder_17bit_yjy # (.UUID(64'd4190818314632917732 ^ UUID)) adder_17bit_yjy_16 (.clk(clk), .rst(rst), .Input_1(wire_41), .Input_2(wire_17), .\17input_1 (wire_24), .\17input_2 (wire_11), .Input_3(1'd0), .\16_sum (wire_49), .\17sum (wire_31), .\17carry ());
  TC_Splitter16 # (.UUID(64'd1233116171020472415 ^ UUID)) Splitter16_17 (.in(wire_4), .out0(wire_5), .out1(wire_10));
  TC_Splitter8 # (.UUID(64'd635017708745103008 ^ UUID)) Splitter8_18 (.in(wire_5), .out0(wire_39), .out1(wire_36), .out2(wire_43), .out3(wire_27), .out4(wire_68), .out5(wire_47), .out6(wire_66), .out7(wire_55));
  TC_Splitter8 # (.UUID(64'd1808923532811563076 ^ UUID)) Splitter8_19 (.in(wire_10), .out0(wire_65), .out1(wire_6), .out2(wire_25), .out3(wire_56), .out4(wire_16), .out5(wire_51), .out6(wire_23), .out7(wire_24));
  TC_Maker16 # (.UUID(64'd3939790085376568009 ^ UUID)) Maker16_20 (.in0(wire_58), .in1(wire_48), .out(wire_41));
  TC_Maker8 # (.UUID(64'd400372928953692755 ^ UUID)) Maker8_21 (.in0(1'd0), .in1(wire_39), .in2(wire_36), .in3(wire_43), .in4(wire_27), .in5(wire_68), .in6(wire_47), .in7(wire_66), .out(wire_58));
  TC_Maker8 # (.UUID(64'd3003221394930974192 ^ UUID)) Maker8_22 (.in0(wire_55), .in1(wire_65), .in2(wire_6), .in3(wire_25), .in4(wire_56), .in5(wire_16), .in6(wire_51), .in7(wire_23), .out(wire_48));
  TC_Splitter16 # (.UUID(64'd2083224792525235346 ^ UUID)) Splitter16_23 (.in(wire_49), .out0(wire_7), .out1(wire_32));
  TC_Register # (.UUID(64'd221619061319804776 ^ UUID), .BIT_WIDTH(64'd8)) Register8_24 (.clk(clk), .rst(rst), .load(wire_15), .save(wire_13), .in(wire_1), .out(wire_22));
  TC_Register # (.UUID(64'd2610169882889075233 ^ UUID), .BIT_WIDTH(64'd8)) Register8_25 (.clk(clk), .rst(rst), .load(wire_15), .save(wire_13), .in(wire_30), .out(wire_45));
  TC_Mux # (.UUID(64'd1680111872412221545 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_26 (.sel(wire_2), .in0(wire_7), .in1(8'd0), .out(wire_1));
  TC_Mux # (.UUID(64'd2496844361308527249 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_27 (.sel(wire_2), .in0(wire_32), .in1(8'd0), .out(wire_30));
  TC_Mux # (.UUID(64'd1658352251236552184 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_28 (.sel(wire_13), .in0(wire_22), .in1(wire_1), .out(wire_37));
  TC_Mux # (.UUID(64'd2249757272663880783 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_29 (.sel(wire_13), .in0(wire_45), .in1(wire_30), .out(wire_62));
  TC_Not # (.UUID(64'd926199163605819017 ^ UUID), .BIT_WIDTH(64'd1)) Not_30 (.in(wire_13), .out(wire_15));
  TC_Register # (.UUID(64'd2021916122347157632 ^ UUID), .BIT_WIDTH(64'd8)) Register8_31 (.clk(clk), .rst(rst), .load(wire_15), .save(wire_13), .in(wire_35), .out(wire_67));
  TC_Mux # (.UUID(64'd3054031882490479354 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_32 (.sel(wire_2), .in0({{7{1'b0}}, wire_31 }), .in1(8'd0), .out(wire_35));
  TC_Mux # (.UUID(64'd3404426579113265709 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_33 (.sel(wire_13), .in0(wire_67), .in1(wire_35), .out(wire_26));

  wire [15:0] wire_0;
  wire [7:0] wire_1;
  wire [0:0] wire_2;
  wire [0:0] wire_3;
  wire [15:0] wire_4;
  wire [7:0] wire_5;
  wire [0:0] wire_6;
  wire [7:0] wire_7;
  wire [7:0] wire_8;
  wire [7:0] wire_9;
  wire [7:0] wire_10;
  wire [0:0] wire_11;
  wire [63:0] wire_12;
  assign wire_12 = i_msg_64;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  assign wire_14 = clk;
  wire [0:0] wire_15;
  wire [0:0] wire_16;
  wire [15:0] wire_17;
  wire [31:0] wire_18;
  wire [63:0] wire_19;
  wire [15:0] wire_20;
  wire [63:0] wire_21;
  wire [7:0] wire_22;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  wire [7:0] wire_26;
  assign Output_1 = wire_26;
  wire [0:0] wire_27;
  wire [63:0] wire_28;
  wire [7:0] wire_29;
  wire [7:0] wire_30;
  wire [0:0] wire_31;
  wire [7:0] wire_32;
  wire [7:0] wire_33;
  wire [7:0] wire_34;
  wire [7:0] wire_35;
  wire [0:0] wire_36;
  wire [7:0] wire_37;
  assign Output_2 = wire_37;
  wire [7:0] wire_38;
  wire [0:0] wire_39;
  wire [7:0] wire_40;
  wire [15:0] wire_41;
  wire [31:0] wire_42;
  wire [0:0] wire_43;
  wire [15:0] wire_44;
  wire [7:0] wire_45;
  wire [7:0] wire_46;
  wire [0:0] wire_47;
  wire [7:0] wire_48;
  wire [15:0] wire_49;
  wire [7:0] wire_50;
  wire [0:0] wire_51;
  wire [7:0] wire_52;
  wire [15:0] wire_53;
  wire [7:0] wire_54;
  wire [0:0] wire_55;
  wire [0:0] wire_56;
  wire [7:0] wire_57;
  wire [7:0] wire_58;
  wire [7:0] wire_59;
  wire [7:0] wire_60;
  wire [7:0] wire_61;
  wire [7:0] wire_62;
  assign Output_3 = wire_62;
  wire [0:0] wire_63;
  assign wire_63 = rstn;
  wire [7:0] wire_64;
  wire [0:0] wire_65;
  wire [0:0] wire_66;
  wire [7:0] wire_67;
  wire [0:0] wire_68;

endmodule
