module mulMiddle_4_2_yjy (clk, rst, clk, rstn, i_msg_64, Output_1, Output_2);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [0:0] clk;
  input  wire [0:0] rstn;
  input  wire [63:0] i_msg_64;
  output  wire [7:0] Output_1;
  output  wire [15:0] Output_2;

  TC_Register # (.UUID(64'd3335127615014970555 ^ UUID), .BIT_WIDTH(64'd64)) Register64_0 (.clk(clk), .rst(rst), .load(wire_9), .save(wire_8), .in(wire_1), .out(wire_0));
  TC_Not # (.UUID(64'd2531310591324011899 ^ UUID), .BIT_WIDTH(64'd1)) Not_1 (.in(wire_44), .out(wire_2));
  TC_Or # (.UUID(64'd3621129731518956724 ^ UUID), .BIT_WIDTH(64'd1)) Or_2 (.in0(wire_62), .in1(wire_2), .out(wire_8));
  TC_Not # (.UUID(64'd597646915276082570 ^ UUID), .BIT_WIDTH(64'd1)) Not_3 (.in(wire_8), .out(wire_9));
  TC_Mux # (.UUID(64'd3795879347822337203 ^ UUID), .BIT_WIDTH(64'd64)) Mux64_4 (.sel(wire_2), .in0(wire_3), .in1(64'd0), .out(wire_1));
  TC_Mux # (.UUID(64'd696410714065915029 ^ UUID), .BIT_WIDTH(64'd64)) Mux64_5 (.sel(wire_8), .in0(wire_0), .in1(wire_1), .out(wire_46));
  TC_Splitter64 # (.UUID(64'd1543269868205825844 ^ UUID)) Splitter64_6 (.in(wire_46), .out0(wire_21), .out1(wire_38), .out2(wire_34), .out3(wire_37), .out4(wire_16), .out5(wire_45), .out6(wire_32), .out7(wire_30));
  TC_Maker32 # (.UUID(64'd1403451493815708811 ^ UUID)) Maker32_7 (.in0(wire_21), .in1(wire_38), .in2(wire_34), .in3(wire_37), .out(wire_50));
  TC_Maker32 # (.UUID(64'd3899840429335718740 ^ UUID)) Maker32_8 (.in0(wire_16), .in1(wire_45), .in2(wire_32), .in3(wire_30), .out(wire_52));
  TC_Splitter32 # (.UUID(64'd1592713307114091917 ^ UUID)) Splitter32_9 (.in(wire_50), .out0(wire_43), .out1(wire_56), .out2(wire_18), .out3());
  TC_Splitter32 # (.UUID(64'd4244626464549385563 ^ UUID)) Splitter32_10 (.in(wire_52), .out0(wire_60), .out1(wire_6), .out2(wire_4), .out3());
  TC_Splitter16 # (.UUID(64'd3278721336715845588 ^ UUID)) Splitter16_11 (.in(wire_11), .out0(wire_39), .out1(wire_61));
  TC_Splitter8 # (.UUID(64'd3398467665959443233 ^ UUID)) Splitter8_12 (.in(wire_39), .out0(wire_53), .out1(wire_24), .out2(wire_67), .out3(wire_13), .out4(wire_58), .out5(wire_48), .out6(wire_7), .out7(wire_26));
  TC_Splitter8 # (.UUID(64'd3094421939014464040 ^ UUID)) Splitter8_13 (.in(wire_61), .out0(wire_55), .out1(wire_54), .out2(wire_42), .out3(wire_40), .out4(wire_22), .out5(wire_23), .out6(wire_19), .out7(wire_49));
  TC_Maker16 # (.UUID(64'd4223464890521494382 ^ UUID)) Maker16_14 (.in0(wire_65), .in1(wire_15), .out(wire_63));
  TC_Maker8 # (.UUID(64'd1737968322881990338 ^ UUID)) Maker8_15 (.in0(1'd0), .in1(wire_53), .in2(wire_24), .in3(wire_67), .in4(wire_13), .in5(wire_58), .in6(wire_48), .in7(wire_7), .out(wire_65));
  TC_Maker8 # (.UUID(64'd547079170662861938 ^ UUID)) Maker8_16 (.in0(wire_26), .in1(wire_55), .in2(wire_54), .in3(wire_42), .in4(wire_40), .in5(wire_22), .in6(wire_23), .in7(wire_19), .out(wire_15));
  TC_Splitter16 # (.UUID(64'd338397297918324923 ^ UUID)) Splitter16_17 (.in(wire_10), .out0(wire_51), .out1(wire_36));
  TC_Register # (.UUID(64'd452998064826846838 ^ UUID), .BIT_WIDTH(64'd8)) Register8_18 (.clk(clk), .rst(rst), .load(wire_25), .save(wire_8), .in(wire_17), .out(wire_41));
  TC_Register # (.UUID(64'd3043137702760234011 ^ UUID), .BIT_WIDTH(64'd8)) Register8_19 (.clk(clk), .rst(rst), .load(wire_25), .save(wire_8), .in(wire_5), .out(wire_29));
  TC_Mux # (.UUID(64'd4599645262819705720 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_20 (.sel(wire_2), .in0(wire_51), .in1(8'd0), .out(wire_17));
  TC_Mux # (.UUID(64'd1103413142931993449 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_21 (.sel(wire_2), .in0(wire_36), .in1(8'd0), .out(wire_5));
  TC_Mux # (.UUID(64'd1389974664402648354 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_22 (.sel(wire_8), .in0(wire_41), .in1(wire_17), .out(wire_47));
  TC_Mux # (.UUID(64'd285418302731830080 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_23 (.sel(wire_8), .in0(wire_29), .in1(wire_5), .out(wire_57));
  TC_Not # (.UUID(64'd1375626209822625454 ^ UUID), .BIT_WIDTH(64'd1)) Not_24 (.in(wire_8), .out(wire_25));
  TC_Register # (.UUID(64'd2026819161103719471 ^ UUID), .BIT_WIDTH(64'd8)) Register8_25 (.clk(clk), .rst(rst), .load(wire_25), .save(wire_8), .in(wire_31), .out(wire_33));
  TC_Mux # (.UUID(64'd427053304534288437 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_26 (.sel(wire_2), .in0({{7{1'b0}}, wire_35 }), .in1(8'd0), .out(wire_31));
  TC_Mux # (.UUID(64'd4103048019201211416 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_27 (.sel(wire_8), .in0(wire_33), .in1(wire_31), .out(wire_66));
  mul8_top_yjy # (.UUID(64'd2584806280345030785 ^ UUID)) mul8_top_yjy_28 (.clk(clk), .rst(rst), .wi_a_8bit(wire_43), .wi_b_8bit(wire_4), .Output(wire_59));
  mul8_top_yjy # (.UUID(64'd3244768142473780112 ^ UUID)) mul8_top_yjy_29 (.clk(clk), .rst(rst), .wi_a_8bit(wire_56), .wi_b_8bit(wire_6), .Output(wire_64));
  mul8_top_yjy # (.UUID(64'd4038594491351837280 ^ UUID)) mul8_top_yjy_30 (.clk(clk), .rst(rst), .wi_a_8bit(wire_18), .wi_b_8bit(wire_60), .Output(wire_28));
  mul8_top_yjy # (.UUID(64'd1546624918859298927 ^ UUID)) mul8_top_yjy_31 (.clk(clk), .rst(rst), .wi_a_8bit(8'd0), .wi_b_8bit(8'd0), .Output(wire_14));
  Compr42with16Bits_yjy # (.UUID(64'd237150703604327293 ^ UUID)) Compr42with16Bits_yjy_32 (.clk(clk), .rst(rst), .Input_1(wire_59), .Input_2(wire_64), .Input_3(wire_28), .Input_4(wire_14), .\1_out (wire_20), .sum(wire_12), .carr(wire_11));
  adder_17bit_yjy # (.UUID(64'd2657036286860137600 ^ UUID)) adder_17bit_yjy_33 (.clk(clk), .rst(rst), .Input_1(wire_63), .Input_2(wire_12), .\17input_1 (wire_49), .\17input_2 (wire_20), .Input_3(1'd0), .\16_sum (wire_10), .\17sum (wire_35), .\17carry ());
  TC_Maker16 # (.UUID(64'd2380114090928370134 ^ UUID)) Maker16_34 (.in0(wire_47), .in1(wire_57), .out(wire_27));

  wire [63:0] wire_0;
  wire [63:0] wire_1;
  wire [0:0] wire_2;
  wire [63:0] wire_3;
  assign wire_3 = i_msg_64;
  wire [7:0] wire_4;
  wire [7:0] wire_5;
  wire [7:0] wire_6;
  wire [0:0] wire_7;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  wire [15:0] wire_10;
  wire [15:0] wire_11;
  wire [15:0] wire_12;
  wire [0:0] wire_13;
  wire [15:0] wire_14;
  wire [7:0] wire_15;
  wire [7:0] wire_16;
  wire [7:0] wire_17;
  wire [7:0] wire_18;
  wire [0:0] wire_19;
  wire [0:0] wire_20;
  wire [7:0] wire_21;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [15:0] wire_27;
  assign Output_2 = wire_27;
  wire [15:0] wire_28;
  wire [7:0] wire_29;
  wire [7:0] wire_30;
  wire [7:0] wire_31;
  wire [7:0] wire_32;
  wire [7:0] wire_33;
  wire [7:0] wire_34;
  wire [0:0] wire_35;
  wire [7:0] wire_36;
  wire [7:0] wire_37;
  wire [7:0] wire_38;
  wire [7:0] wire_39;
  wire [0:0] wire_40;
  wire [7:0] wire_41;
  wire [0:0] wire_42;
  wire [7:0] wire_43;
  wire [0:0] wire_44;
  assign wire_44 = rstn;
  wire [7:0] wire_45;
  wire [63:0] wire_46;
  wire [7:0] wire_47;
  wire [0:0] wire_48;
  wire [0:0] wire_49;
  wire [31:0] wire_50;
  wire [7:0] wire_51;
  wire [31:0] wire_52;
  wire [0:0] wire_53;
  wire [0:0] wire_54;
  wire [0:0] wire_55;
  wire [7:0] wire_56;
  wire [7:0] wire_57;
  wire [0:0] wire_58;
  wire [15:0] wire_59;
  wire [7:0] wire_60;
  wire [7:0] wire_61;
  wire [0:0] wire_62;
  assign wire_62 = clk;
  wire [15:0] wire_63;
  wire [15:0] wire_64;
  wire [7:0] wire_65;
  wire [7:0] wire_66;
  assign Output_1 = wire_66;
  wire [0:0] wire_67;

endmodule
