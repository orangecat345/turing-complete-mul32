module mul_top_yjy (clk, rst, clk, i_msg, rstn, delay_4, Output_1, Output_2, Output_3, high_result);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [0:0] clk;
  input  wire [63:0] i_msg;
  input  wire [0:0] rstn;
  output  wire [0:0] delay_4;
  output  wire [31:0] Output_1;
  output  wire [31:0] Output_2;
  output  wire [31:0] Output_3;
  output  wire [31:0] high_result;

  TC_Maker32 # (.UUID(64'd491013554895460409 ^ UUID)) Maker32_0 (.in0(8'd0), .in1(wire_50), .in2(wire_14), .in3(wire_53), .out(wire_19));
  TC_Splitter16 # (.UUID(64'd1178369419794067826 ^ UUID)) Splitter16_1 (.in(wire_9), .out0(wire_50), .out1(wire_14));
  TC_Maker32 # (.UUID(64'd3790761036020857293 ^ UUID)) Maker32_2 (.in0(wire_20), .in1(wire_3), .in2(wire_58), .in3(wire_45), .out(wire_15));
  TC_Splitter16 # (.UUID(64'd152569839927454265 ^ UUID)) Splitter16_3 (.in(wire_49), .out0(wire_20), .out1(wire_3));
  TC_Splitter16 # (.UUID(64'd4141198415988714931 ^ UUID)) Splitter16_4 (.in(wire_5), .out0(wire_58), .out1(wire_45));
  TC_Maker32 # (.UUID(64'd632314921896204275 ^ UUID)) Maker32_5 (.in0(wire_44), .in1(wire_28), .in2(wire_32), .in3(wire_55), .out(wire_36));
  TC_Splitter16 # (.UUID(64'd4050665473848537250 ^ UUID)) Splitter16_6 (.in(wire_43), .out0(wire_28), .out1(wire_32));
  TC_Maker32 # (.UUID(64'd2812620014313922675 ^ UUID)) Maker32_7 (.in0(wire_12), .in1(wire_24), .in2(wire_57), .in3(wire_23), .out(wire_48));
  TC_Splitter16 # (.UUID(64'd3631752085026053919 ^ UUID)) Splitter16_8 (.in(wire_25), .out0(wire_57), .out1(wire_23));
  TC_Splitter16 # (.UUID(64'd2890889190553753470 ^ UUID)) Splitter16_9 (.in(wire_33), .out0(wire_12), .out1(wire_24));
  TC_Maker32 # (.UUID(64'd507656039066428653 ^ UUID)) Maker32_10 (.in0(wire_11), .in1(wire_16), .in2(wire_46), .in3(8'd0), .out(wire_27));
  TC_Mul # (.UUID(64'd2691410044601611021 ^ UUID), .BIT_WIDTH(64'd32)) Mul32_11 (.in0(wire_8), .in1(wire_17), .out0(wire_22), .out1(wire_21));
  TC_Splitter64 # (.UUID(64'd2500474701101987968 ^ UUID)) Splitter64_12 (.in(wire_0), .out0(wire_51), .out1(wire_4), .out2(wire_29), .out3(wire_40), .out4(wire_35), .out5(wire_54), .out6(wire_56), .out7(wire_6));
  TC_Maker32 # (.UUID(64'd3315045708623855349 ^ UUID)) Maker32_13 (.in0(wire_51), .in1(wire_4), .in2(wire_29), .in3(wire_40), .out(wire_8));
  TC_Maker32 # (.UUID(64'd640275572284684509 ^ UUID)) Maker32_14 (.in0(wire_35), .in1(wire_54), .in2(wire_56), .in3(wire_6), .out(wire_17));
  TC_Constant # (.UUID(64'd1372811850642340322 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_15 (.out(wire_10));
  TC_Not # (.UUID(64'd4246925385856427608 ^ UUID), .BIT_WIDTH(64'd1)) Not_16 (.in(wire_52), .out(wire_26));
  TC_DelayLine # (.UUID(64'd2962909952648258708 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_17 (.clk(clk), .rst(rst), .in(wire_1), .out(wire_47));
  TC_DelayLine # (.UUID(64'd298069981974059390 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_18 (.clk(clk), .rst(rst), .in(wire_47), .out(wire_7));
  TC_DelayLine # (.UUID(64'd2736359972295435874 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_19 (.clk(clk), .rst(rst), .in(wire_7), .out(wire_34));
  TC_Or3 # (.UUID(64'd2082453249592269091 ^ UUID), .BIT_WIDTH(64'd1)) Or3_20 (.in0(wire_34), .in1(1'd0), .in2(1'd0), .out(wire_39));
  mulMiddle_4_1_yjy # (.UUID(64'd882715702263392216 ^ UUID)) mulMiddle_4_1_yjy_21 (.clk(clk), .rst(rst), .clk(wire_1), .rstn(wire_10), .i_msg_64(wire_0), .Output_1(wire_16), .Output_2(wire_18), .Output_3(wire_44));
  mult_8_1_8bit_hso # (.UUID(64'd1868010957065212696 ^ UUID)) mult_8_1_8bit_hso_22 (.clk(clk), .rst(rst), .i_msg_64(wire_0), .clk(wire_1), .rstn(wire_10), .low_result_16bit(wire_49));
  adder_8bit_yjy # (.UUID(64'd3415230542068637573 ^ UUID)) adder_8bit_yjy_23 (.clk(clk), .rst(rst), .Input_1(wire_18), .Input_2(wire_2), .Input_3(1'd0), .Output_1(wire_53), .Output_2(wire_42));
  adder_32bit_lgy # (.UUID(64'd1244611914891560576 ^ UUID)) adder_32bit_lgy_24 (.clk(clk), .rst(rst), .Input_1(wire_19), .Input_2(wire_15), .Input_3(1'd0), .rstn(wire_10), .clk(wire_1), .Output_1(wire_31), .Output_2(wire_38));
  adder_8bit_yjy # (.UUID(64'd3887797524087931119 ^ UUID)) adder_8bit_yjy_25 (.clk(clk), .rst(rst), .Input_1(wire_37), .Input_2(wire_42), .Input_3(1'd0), .Output_1(wire_30), .Output_2());
  adder_8bit_yjy # (.UUID(64'd2160155339316910245 ^ UUID)) adder_8bit_yjy_26 (.clk(clk), .rst(rst), .Input_1(wire_30), .Input_2(wire_38), .Input_3(1'd0), .Output_1(wire_11), .Output_2());
  mulMiddle_4_2_yjy # (.UUID(64'd318064441174018236 ^ UUID)) mulMiddle_4_2_yjy_27 (.clk(clk), .rst(rst), .clk(wire_1), .rstn(wire_10), .i_msg_64(wire_0), .Output_1(wire_37), .Output_2(wire_5));
  mulMiddle_4_3_yjy # (.UUID(64'd4053004592916859895 ^ UUID)) mulMiddle_4_3_yjy_28 (.clk(clk), .rst(rst), .clk(wire_1), .rstn(wire_10), .i_msg_64(wire_0), .Output_1(wire_46), .Output_2(wire_33));
  mulMiddle_2_2_yjy # (.UUID(64'd1671485050718566416 ^ UUID)) mulMiddle_2_2_yjy_29 (.clk(clk), .rst(rst), .clk(wire_1), .rstn(wire_10), .Input(wire_0), .Output_1(wire_55), .Output_2(wire_43));
  mult_8_2_8bit_hso # (.UUID(64'd3625949718049989348 ^ UUID)) mult_8_2_8bit_hso_30 (.clk(clk), .rst(rst), .i_msg_64(wire_0), .clk(wire_1), .rstn(wire_10), .low_result_16bit(wire_25));
  adder_32bit_lgy # (.UUID(64'd1700948130532912039 ^ UUID)) adder_32bit_lgy_31 (.clk(clk), .rst(rst), .Input_1(wire_13), .Input_2(wire_27), .Input_3(1'd0), .rstn(wire_10), .clk(wire_1), .Output_1(wire_41), .Output_2());
  adder_32bit_lgy # (.UUID(64'd1837899594163424462 ^ UUID)) adder_32bit_lgy_32 (.clk(clk), .rst(rst), .Input_1(wire_36), .Input_2(wire_48), .Input_3(1'd0), .rstn(wire_10), .clk(wire_1), .Output_1(wire_13), .Output_2());
  mulMiddle_2_1_yjy # (.UUID(64'd2775608885769112211 ^ UUID)) mulMiddle_2_1_yjy_33 (.clk(clk), .rst(rst), .clk(wire_1), .rstn(wire_10), .Input(wire_0), .Output_1(wire_2), .Output_2(wire_9));

  wire [63:0] wire_0;
  assign wire_0 = i_msg;
  wire [0:0] wire_1;
  assign wire_1 = clk;
  wire [7:0] wire_2;
  wire [7:0] wire_3;
  wire [7:0] wire_4;
  wire [15:0] wire_5;
  wire [7:0] wire_6;
  wire [0:0] wire_7;
  wire [31:0] wire_8;
  wire [15:0] wire_9;
  wire [0:0] wire_10;
  wire [7:0] wire_11;
  wire [7:0] wire_12;
  wire [31:0] wire_13;
  wire [7:0] wire_14;
  wire [31:0] wire_15;
  wire [7:0] wire_16;
  wire [31:0] wire_17;
  wire [7:0] wire_18;
  wire [31:0] wire_19;
  wire [7:0] wire_20;
  wire [31:0] wire_21;
  assign Output_2 = wire_21;
  wire [31:0] wire_22;
  assign Output_1 = wire_22;
  wire [7:0] wire_23;
  wire [7:0] wire_24;
  wire [15:0] wire_25;
  wire [0:0] wire_26;
  wire [31:0] wire_27;
  wire [7:0] wire_28;
  wire [7:0] wire_29;
  wire [7:0] wire_30;
  wire [31:0] wire_31;
  assign Output_3 = wire_31;
  wire [7:0] wire_32;
  wire [15:0] wire_33;
  wire [0:0] wire_34;
  wire [7:0] wire_35;
  wire [31:0] wire_36;
  wire [7:0] wire_37;
  wire [7:0] wire_38;
  wire [0:0] wire_39;
  assign delay_4 = wire_39;
  wire [7:0] wire_40;
  wire [31:0] wire_41;
  assign high_result = wire_41;
  wire [7:0] wire_42;
  wire [15:0] wire_43;
  wire [7:0] wire_44;
  wire [7:0] wire_45;
  wire [7:0] wire_46;
  wire [0:0] wire_47;
  wire [31:0] wire_48;
  wire [15:0] wire_49;
  wire [7:0] wire_50;
  wire [7:0] wire_51;
  wire [0:0] wire_52;
  assign wire_52 = 0;
  wire [7:0] wire_53;
  wire [7:0] wire_54;
  wire [7:0] wire_55;
  wire [7:0] wire_56;
  wire [7:0] wire_57;
  wire [7:0] wire_58;

endmodule
